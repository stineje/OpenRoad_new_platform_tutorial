A behavioral module for both a CLKGATE and LATCH need to be included in the platforms directory and their respective paths added into the config.mk file. Refer to another platform to get an idea on how these are constructed.
